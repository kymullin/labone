/*-------------------------------------------------------------
    Project Lab 1 - Main Project
       Program by: Zachary Bonneau
    Creation Date: 
     Program Name: 
    SubProgram of: 
  
    Program Description:
    

    Inputs:
        
    
    Outputs:
       

*///-----------------------------------------------------------

// directive calls


// module code here
module <name>(

);


endmodule